// ---------------------------------------------------------------------------------------
// File               : gen_top_asrt_if.sv
// Version            : 
// Author             : 
// ---------------------------------------------------------------------------------------
// Description        : Generated assertion interface binded to the
//                      top module
// ---------------------------------------------------------------------------------------


// =======================================================================================
//  Interface:       top_asrt_if
// ---------------------------------------------------------------------------------------
//
//  Generated assertion interface. Binded to the top DUT from the testbench.
//  Includes variables, models, properties, and assertions.
//
//  Parameters:
//    WIDTH
//
//  Ports:
//    clk
//    rst
//    data_in
//    data_out
//    ctrl
//
// =======================================================================================

interface top_asrt_if #( 
    parameter logic [3:0] WIDTH = 8  
) (
  input logic              clk,
  input logic              rst,
  input logic [WIDTH-1:0]  data_in,
  input logic [WIDTH-1:0]  data_out,
  input keys_s             ctrl
);

  // =====================================================================================
  //                                                                            Data Types
  // =====================================================================================

  // =====================================================================================
  //                                                                            Parameters
  // =====================================================================================

  `define PATH_TOP  = i_dut

  // =====================================================================================
  //                                                                    Imports & Includes
  // =====================================================================================

  // =====================================================================================
  //                                                                             Variables
  // =====================================================================================

  //---------------------------------------PORTS----------------------------------------//

  //----------------------------------------FIFO----------------------------------------//

  // var: i_rx_i_fifo_data_out
  logic [WIDTH-1 : 0]                 i_rx_i_fifo_data_out;

  //-----------------------------------------TX-----------------------------------------//

  // var: txd
  logic                               txd;

  //-----------------------------------------RX-----------------------------------------//

  // var: rxd
  logic                               rxd;

  //----------------------------------------FIFO----------------------------------------//

  // var: re
  logic                               re;

  // var: we
  logic                               we;

  //-------------------------------------REGISTERS--------------------------------------//

  //----------------------------------------TOP-----------------------------------------//

  // var: addr_s
  logic [1:0]                         addr_s;

  // var: laddr_s
  logic [c_VERY_LOOONG_ADDR - 1 : 0]  laddr_s;

  // var: start_s
  logic                               start_s;

  // var: we_s
  logic                               we_s;

  // var: data_s
  data_t                              data_s;

  //-----------------------------------------TX-----------------------------------------//

  // var: tx_s
  logic                               tx_s;

  //-----------------------------------------RX-----------------------------------------//

  // var: rx_s
  logic                               rx_s;

  //----------------------------------------FIFO----------------------------------------//

  // var: data_s
  logic [WIDTH-1 : 0]                 data_s;
  
  //----------------------------------Models variables----------------------------------//

  // =====================================================================================
  //                                                                                Models
  // =====================================================================================

  // =====================================================================================
  //                                                                    Output Assignments
  // =====================================================================================

  assign i_rx_i_fifo_data_out = `PATH_TOP.i_rx.i_fifo.data_out;
  assign txd                  = `PATH_TOP.i_tx.txd;
  assign rxd                  = `PATH_TOP.i_rx.rxd;
  assign re                   = `PATH_TOP.i_rx.i_fifo.re;
  assign we                   = `PATH_TOP.i_rx.i_fifo.we;
  assign addr_s               = `PATH_TOP.addr_s;
  assign laddr_s              = `PATH_TOP.laddr_s;
  assign start_s              = `PATH_TOP.start_s;
  assign we_s                 = `PATH_TOP.we_s;
  assign data_s               = `PATH_TOP.data_s;
  assign tx_s                 = `PATH_TOP.i_tx.tx_s;
  assign rx_s                 = `PATH_TOP.i_rx.rx_s;
  assign data_s               = `PATH_TOP.i_rx.i_fifo.data_s;

  // =====================================================================================
  //                                                                     Common Properties
  // =====================================================================================

  //                ______________
  // SIG: _________/  \___________
  //             __
  // COND: _____/  \______________
  property COND_ROSE_ACTIVE_SIGNAL_NEXT_CYCLE(COND, SIG);
    $rose(COND) |=> SIG;
  endproperty
    
  // =====================================================================================
  //                                                                            Assertions
  // =====================================================================================
  // `include "assertions_include_file_example.svh"

endinterface : top_asrt_if

// =======================================================================================
//                                                                             End-Of-File
// =======================================================================================