module tx #(
    parameter logic [3:0] WIDTH = 8  
)(
    input logic clk,
    input logic rst,
    output logic txd
);
  logic tx_c, tx_s;
  
endmodule